module ControlUnit(opcode,funct);
    input [5:0] opcode;
    input [5:0] funct;
endmodule